//////////////////////////////
// һά����Ҷ�任��֤ƽ̨����
//////////////////////////////

`timescale 1ns/1ps
module fft_matrix_tb(
    
);

